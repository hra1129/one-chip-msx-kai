module tb;
	localparam		CLK_BASE	= 1000000000/21480;

	reg					CLK21M;
	reg					RESET;
	reg			[ 1:0]	DOTSTATE;
	reg			[ 2:0]	EIGHTDOTSTATE;
	reg			[ 8:0]	DOTCOUNTERX;
	reg			[ 8:0]	DOTCOUNTERYP;
	reg					BWINDOW_Y;
	wire				PVDPS0SPCOLLISIONINCIDENCE;
	wire				PVDPS0SPOVERMAPPED;
	wire		[ 4:0]	PVDPS0SPOVERMAPPEDNUM;
	wire		[ 8:0]	PVDPS3S4SPCOLLISIONX;
	wire		[ 8:0]	PVDPS5S6SPCOLLISIONY;
	reg					PVDPS0RESETREQ;
	wire				PVDPS0RESETACK;
	reg					PVDPS5RESETREQ;
	wire				PVDPS5RESETACK;
	reg					REG_R1_SP_SIZE;
	reg					REG_R1_SP_ZOOM;
	reg			[ 9:0]	REG_R11R5_SP_ATR_ADDR;
	reg			[ 5:0]	REG_R6_SP_GEN_ADDR;
	reg					REG_R8_COL0_ON;
	reg					REG_R8_SP_OFF;
	reg			[ 7:0]	REG_R23_VSTART_LINE;
	reg			[ 2:0]	REG_R27_H_SCROLL;
	reg					SPMODE2;
	reg					VRAMINTERLEAVEMODE;
	wire				SPVRAMACCESSING;
	reg			[ 7:0]	PRAMDAT;
	wire		[16:0]	PRAMADR;
	wire				SPCOLOROUT;
	wire		[ 3:0]	SPCOLORCODE;

	reg			[ 7:0]	virtual_vram[longint unsigned];
	integer				vram_address;

	// -------------------------------------------------------------
	//	clock generator
	// -------------------------------------------------------------
	always #(CLK_BASE/2) begin
		CLK21M	<= ~CLK21M;
	end

	// -------------------------------------------------------------
	//	DUT
	// -------------------------------------------------------------
	VDP_SPRITE u_dut (
		.CLK21M							( CLK21M						),
		.RESET							( RESET							),
		.DOTSTATE						( DOTSTATE						),
		.EIGHTDOTSTATE					( EIGHTDOTSTATE					),
		.DOTCOUNTERX					( DOTCOUNTERX					),
		.DOTCOUNTERYP					( DOTCOUNTERYP					),
		.BWINDOW_Y						( BWINDOW_Y						),
		.PVDPS0SPCOLLISIONINCIDENCE		( PVDPS0SPCOLLISIONINCIDENCE	),
		.PVDPS0SPOVERMAPPED				( PVDPS0SPOVERMAPPED			),
		.PVDPS0SPOVERMAPPEDNUM			( PVDPS0SPOVERMAPPEDNUM			),
		.PVDPS3S4SPCOLLISIONX			( PVDPS3S4SPCOLLISIONX			),
		.PVDPS5S6SPCOLLISIONY			( PVDPS5S6SPCOLLISIONY			),
		.PVDPS0RESETREQ					( PVDPS0RESETREQ				),
		.PVDPS0RESETACK					( PVDPS0RESETACK				),
		.PVDPS5RESETREQ					( PVDPS5RESETREQ				),
		.PVDPS5RESETACK					( PVDPS5RESETACK				),
		.REG_R1_SP_SIZE					( REG_R1_SP_SIZE				),
		.REG_R1_SP_ZOOM					( REG_R1_SP_ZOOM				),
		.REG_R11R5_SP_ATR_ADDR			( REG_R11R5_SP_ATR_ADDR			),
		.REG_R6_SP_GEN_ADDR				( REG_R6_SP_GEN_ADDR			),
		.REG_R8_COL0_ON					( REG_R8_COL0_ON				),
		.REG_R8_SP_OFF					( REG_R8_SP_OFF					),
		.REG_R23_VSTART_LINE			( REG_R23_VSTART_LINE			),
		.REG_R27_H_SCROLL				( REG_R27_H_SCROLL				),
		.SPMODE2						( SPMODE2						),
		.VRAMINTERLEAVEMODE				( VRAMINTERLEAVEMODE			),
		.SPVRAMACCESSING				( SPVRAMACCESSING				),
		.PRAMDAT						( PRAMDAT						),
		.PRAMADR						( PRAMADR						),
		.SPCOLOROUT						( SPCOLOROUT					),
		.SPCOLORCODE					( SPCOLORCODE					)
	);

	always @( posedge RESET or posedge CLK21M ) begin
		if( RESET ) begin
			DOTSTATE	<= 2'b10;
		end
		else begin
			case( DOTSTATE )
			2'b00:		DOTSTATE <= 2'b01;
			2'b01:		DOTSTATE <= 2'b11;
			2'b11:		DOTSTATE <= 2'b10;
			2'b10:		DOTSTATE <= 2'b00;
			default:	DOTSTATE <= 2'b00;
			endcase
		end
	end

	always @( posedge RESET or posedge CLK21M ) begin
		if( RESET ) begin
			EIGHTDOTSTATE	<= 3'd0;
		end
		else if( DOTSTATE == 2'b10 ) begin
			EIGHTDOTSTATE	<= DOTCOUNTERX[2:0];
		end
		else begin
			//	hold
		end
	end

	always @( posedge RESET or posedge CLK21M ) begin
		if( RESET ) begin
			DOTCOUNTERX		<= -9'd8;
		end
		else if( DOTSTATE == 2'b11 ) begin
			if( DOTCOUNTERX == 9'd341 ) begin
				DOTCOUNTERX <= -9'd8;
			end
			else begin
				DOTCOUNTERX <= DOTCOUNTERX + 9'd1;
			end
		end
		else begin
			//	hold
		end
	end

	always @( posedge RESET or posedge CLK21M ) begin
		if( RESET ) begin
			DOTCOUNTERYP		<= -9'd8;
		end
		else if( DOTSTATE == 2'b10 && DOTCOUNTERX == 9'd341 ) begin
			if( DOTCOUNTERYP == 9'd264 ) begin
				DOTCOUNTERYP <= -9'd8;
			end
			else begin
				DOTCOUNTERYP <= DOTCOUNTERYP + 9'd1;
			end
		end
		else begin
			//	hold
		end
	end

	always @( posedge CLK21M ) begin
		vram_address	<= PRAMADR;
		PRAMDAT			<= virtual_vram[ vram_address ];
	end

	initial begin
		CLK21M		= 0;
		RESET		= 1;

		BWINDOW_Y = 0;
		PVDPS0RESETREQ = 0;
		PVDPS5RESETREQ = 0;
		REG_R1_SP_SIZE = 1;
		REG_R1_SP_ZOOM = 0;
		REG_R11R5_SP_ATR_ADDR = 0;
		REG_R6_SP_GEN_ADDR = 0;
		REG_R8_COL0_ON = 0;
		REG_R8_SP_OFF = 0;
		REG_R23_VSTART_LINE = 0;
		REG_R27_H_SCROLL = 0;
		SPMODE2 = 1;
		VRAMINTERLEAVEMODE = 0;

		virtual_vram[ 17'h07400 ]	= 'h24;
		virtual_vram[ 17'h07401 ]	= 'h24;
		virtual_vram[ 17'h07402 ]	= 'h24;
		virtual_vram[ 17'h07403 ]	= 'h24;
		virtual_vram[ 17'h07404 ]	= 'h24;
		virtual_vram[ 17'h07405 ]	= 'h24;
		virtual_vram[ 17'h07406 ]	= 'h24;
		virtual_vram[ 17'h07407 ]	= 'h24;
		virtual_vram[ 17'h07408 ]	= 'h24;
		virtual_vram[ 17'h07409 ]	= 'h24;
		virtual_vram[ 17'h0740A ]	= 'h24;
		virtual_vram[ 17'h0740B ]	= 'h24;
		virtual_vram[ 17'h0740C ]	= 'h24;
		virtual_vram[ 17'h0740D ]	= 'h24;
		virtual_vram[ 17'h0740E ]	= 'h24;
		virtual_vram[ 17'h0740F ]	= 'h24;
		virtual_vram[ 17'h07410 ]	= 'h24;
		virtual_vram[ 17'h07411 ]	= 'h24;
		virtual_vram[ 17'h07412 ]	= 'h24;
		virtual_vram[ 17'h07413 ]	= 'h24;
		virtual_vram[ 17'h07414 ]	= 'h24;
		virtual_vram[ 17'h07415 ]	= 'h24;
		virtual_vram[ 17'h07416 ]	= 'h24;
		virtual_vram[ 17'h07417 ]	= 'h24;
		virtual_vram[ 17'h07418 ]	= 'h24;
		virtual_vram[ 17'h07419 ]	= 'h24;
		virtual_vram[ 17'h0741A ]	= 'h24;
		virtual_vram[ 17'h0741B ]	= 'h24;
		virtual_vram[ 17'h0741C ]	= 'h24;
		virtual_vram[ 17'h0741D ]	= 'h24;
		virtual_vram[ 17'h0741E ]	= 'h24;
		virtual_vram[ 17'h0741F ]	= 'h24;
		virtual_vram[ 17'h07420 ]	= 'h24;
		virtual_vram[ 17'h07421 ]	= 'h24;
		virtual_vram[ 17'h07422 ]	= 'h24;
		virtual_vram[ 17'h07423 ]	= 'h24;
		virtual_vram[ 17'h07424 ]	= 'h24;
		virtual_vram[ 17'h07425 ]	= 'h24;
		virtual_vram[ 17'h07426 ]	= 'h24;
		virtual_vram[ 17'h07427 ]	= 'h24;
		virtual_vram[ 17'h07428 ]	= 'h24;
		virtual_vram[ 17'h07429 ]	= 'h24;
		virtual_vram[ 17'h0742A ]	= 'h24;
		virtual_vram[ 17'h0742B ]	= 'h24;
		virtual_vram[ 17'h0742C ]	= 'h24;
		virtual_vram[ 17'h0742D ]	= 'h24;
		virtual_vram[ 17'h0742E ]	= 'h24;
		virtual_vram[ 17'h0742F ]	= 'h24;
		virtual_vram[ 17'h07430 ]	= 'h24;
		virtual_vram[ 17'h07431 ]	= 'h24;
		virtual_vram[ 17'h07432 ]	= 'h24;
		virtual_vram[ 17'h07433 ]	= 'h24;
		virtual_vram[ 17'h07434 ]	= 'h24;
		virtual_vram[ 17'h07435 ]	= 'h24;
		virtual_vram[ 17'h07436 ]	= 'h24;
		virtual_vram[ 17'h07437 ]	= 'h24;
		virtual_vram[ 17'h07438 ]	= 'h24;
		virtual_vram[ 17'h07439 ]	= 'h24;
		virtual_vram[ 17'h0743A ]	= 'h24;
		virtual_vram[ 17'h0743B ]	= 'h24;
		virtual_vram[ 17'h0743C ]	= 'h24;
		virtual_vram[ 17'h0743D ]	= 'h24;
		virtual_vram[ 17'h0743E ]	= 'h24;
		virtual_vram[ 17'h0743F ]	= 'h24;
		virtual_vram[ 17'h07440 ]	= 'h24;
		virtual_vram[ 17'h07441 ]	= 'h24;
		virtual_vram[ 17'h07442 ]	= 'h24;
		virtual_vram[ 17'h07443 ]	= 'h24;
		virtual_vram[ 17'h07444 ]	= 'h24;
		virtual_vram[ 17'h07445 ]	= 'h24;
		virtual_vram[ 17'h07446 ]	= 'h24;
		virtual_vram[ 17'h07447 ]	= 'h24;
		virtual_vram[ 17'h07448 ]	= 'h24;
		virtual_vram[ 17'h07449 ]	= 'h24;
		virtual_vram[ 17'h0744A ]	= 'h24;
		virtual_vram[ 17'h0744B ]	= 'h24;
		virtual_vram[ 17'h0744C ]	= 'h24;
		virtual_vram[ 17'h0744D ]	= 'h24;
		virtual_vram[ 17'h0744E ]	= 'h24;
		virtual_vram[ 17'h0744F ]	= 'h24;
		virtual_vram[ 17'h07450 ]	= 'h24;
		virtual_vram[ 17'h07451 ]	= 'h24;
		virtual_vram[ 17'h07452 ]	= 'h24;
		virtual_vram[ 17'h07453 ]	= 'h24;
		virtual_vram[ 17'h07454 ]	= 'h24;
		virtual_vram[ 17'h07455 ]	= 'h24;
		virtual_vram[ 17'h07456 ]	= 'h24;
		virtual_vram[ 17'h07457 ]	= 'h24;
		virtual_vram[ 17'h07458 ]	= 'h24;
		virtual_vram[ 17'h07459 ]	= 'h24;
		virtual_vram[ 17'h0745A ]	= 'h24;
		virtual_vram[ 17'h0745B ]	= 'h24;
		virtual_vram[ 17'h0745C ]	= 'h24;
		virtual_vram[ 17'h0745D ]	= 'h24;
		virtual_vram[ 17'h0745E ]	= 'h24;
		virtual_vram[ 17'h0745F ]	= 'h24;
		virtual_vram[ 17'h07460 ]	= 'h24;
		virtual_vram[ 17'h07461 ]	= 'h24;
		virtual_vram[ 17'h07462 ]	= 'h24;
		virtual_vram[ 17'h07463 ]	= 'h24;
		virtual_vram[ 17'h07464 ]	= 'h24;
		virtual_vram[ 17'h07465 ]	= 'h24;
		virtual_vram[ 17'h07466 ]	= 'h24;
		virtual_vram[ 17'h07467 ]	= 'h24;
		virtual_vram[ 17'h07468 ]	= 'h24;
		virtual_vram[ 17'h07469 ]	= 'h24;
		virtual_vram[ 17'h0746A ]	= 'h24;
		virtual_vram[ 17'h0746B ]	= 'h24;
		virtual_vram[ 17'h0746C ]	= 'h24;
		virtual_vram[ 17'h0746D ]	= 'h24;
		virtual_vram[ 17'h0746E ]	= 'h24;
		virtual_vram[ 17'h0746F ]	= 'h24;
		virtual_vram[ 17'h07470 ]	= 'h24;
		virtual_vram[ 17'h07471 ]	= 'h24;
		virtual_vram[ 17'h07472 ]	= 'h24;
		virtual_vram[ 17'h07473 ]	= 'h24;
		virtual_vram[ 17'h07474 ]	= 'h24;
		virtual_vram[ 17'h07475 ]	= 'h24;
		virtual_vram[ 17'h07476 ]	= 'h24;
		virtual_vram[ 17'h07477 ]	= 'h24;
		virtual_vram[ 17'h07478 ]	= 'h24;
		virtual_vram[ 17'h07479 ]	= 'h24;
		virtual_vram[ 17'h0747A ]	= 'h24;
		virtual_vram[ 17'h0747B ]	= 'h24;
		virtual_vram[ 17'h0747C ]	= 'h24;
		virtual_vram[ 17'h0747D ]	= 'h24;
		virtual_vram[ 17'h0747E ]	= 'h24;
		virtual_vram[ 17'h0747F ]	= 'h24;
		virtual_vram[ 17'h07480 ]	= 'h24;
		virtual_vram[ 17'h07481 ]	= 'h24;
		virtual_vram[ 17'h07482 ]	= 'h24;
		virtual_vram[ 17'h07483 ]	= 'h24;
		virtual_vram[ 17'h07484 ]	= 'h24;
		virtual_vram[ 17'h07485 ]	= 'h24;
		virtual_vram[ 17'h07486 ]	= 'h24;
		virtual_vram[ 17'h07487 ]	= 'h24;
		virtual_vram[ 17'h07488 ]	= 'h24;
		virtual_vram[ 17'h07489 ]	= 'h24;
		virtual_vram[ 17'h0748A ]	= 'h24;
		virtual_vram[ 17'h0748B ]	= 'h24;
		virtual_vram[ 17'h0748C ]	= 'h24;
		virtual_vram[ 17'h0748D ]	= 'h24;
		virtual_vram[ 17'h0748E ]	= 'h24;
		virtual_vram[ 17'h0748F ]	= 'h24;
		virtual_vram[ 17'h07490 ]	= 'h24;
		virtual_vram[ 17'h07491 ]	= 'h24;
		virtual_vram[ 17'h07492 ]	= 'h24;
		virtual_vram[ 17'h07493 ]	= 'h24;
		virtual_vram[ 17'h07494 ]	= 'h24;
		virtual_vram[ 17'h07495 ]	= 'h24;
		virtual_vram[ 17'h07496 ]	= 'h24;
		virtual_vram[ 17'h07497 ]	= 'h24;
		virtual_vram[ 17'h07498 ]	= 'h24;
		virtual_vram[ 17'h07499 ]	= 'h24;
		virtual_vram[ 17'h0749A ]	= 'h24;
		virtual_vram[ 17'h0749B ]	= 'h24;
		virtual_vram[ 17'h0749C ]	= 'h24;
		virtual_vram[ 17'h0749D ]	= 'h24;
		virtual_vram[ 17'h0749E ]	= 'h24;
		virtual_vram[ 17'h0749F ]	= 'h24;
		virtual_vram[ 17'h074A0 ]	= 'h24;
		virtual_vram[ 17'h074A1 ]	= 'h24;
		virtual_vram[ 17'h074A2 ]	= 'h24;
		virtual_vram[ 17'h074A3 ]	= 'h24;
		virtual_vram[ 17'h074A4 ]	= 'h24;
		virtual_vram[ 17'h074A5 ]	= 'h24;
		virtual_vram[ 17'h074A6 ]	= 'h24;
		virtual_vram[ 17'h074A7 ]	= 'h24;
		virtual_vram[ 17'h074A8 ]	= 'h24;
		virtual_vram[ 17'h074A9 ]	= 'h24;
		virtual_vram[ 17'h074AA ]	= 'h24;
		virtual_vram[ 17'h074AB ]	= 'h24;
		virtual_vram[ 17'h074AC ]	= 'h24;
		virtual_vram[ 17'h074AD ]	= 'h24;
		virtual_vram[ 17'h074AE ]	= 'h24;
		virtual_vram[ 17'h074AF ]	= 'h24;
		virtual_vram[ 17'h074B0 ]	= 'h62;
		virtual_vram[ 17'h074B1 ]	= 'h62;
		virtual_vram[ 17'h074B2 ]	= 'h62;
		virtual_vram[ 17'h074B3 ]	= 'h62;
		virtual_vram[ 17'h074B4 ]	= 'h62;
		virtual_vram[ 17'h074B5 ]	= 'h62;
		virtual_vram[ 17'h074B6 ]	= 'h62;
		virtual_vram[ 17'h074B7 ]	= 'h62;
		virtual_vram[ 17'h074B8 ]	= 'h62;
		virtual_vram[ 17'h074B9 ]	= 'h62;
		virtual_vram[ 17'h074BA ]	= 'h62;
		virtual_vram[ 17'h074BB ]	= 'h62;
		virtual_vram[ 17'h074BC ]	= 'h62;
		virtual_vram[ 17'h074BD ]	= 'h62;
		virtual_vram[ 17'h074BE ]	= 'h62;
		virtual_vram[ 17'h074BF ]	= 'h62;
		virtual_vram[ 17'h074C0 ]	= 'h62;
		virtual_vram[ 17'h074C1 ]	= 'h62;
		virtual_vram[ 17'h074C2 ]	= 'h62;
		virtual_vram[ 17'h074C3 ]	= 'h62;
		virtual_vram[ 17'h074C4 ]	= 'h62;
		virtual_vram[ 17'h074C5 ]	= 'h62;
		virtual_vram[ 17'h074C6 ]	= 'h62;
		virtual_vram[ 17'h074C7 ]	= 'h62;
		virtual_vram[ 17'h074C8 ]	= 'h62;
		virtual_vram[ 17'h074C9 ]	= 'h62;
		virtual_vram[ 17'h074CA ]	= 'h62;
		virtual_vram[ 17'h074CB ]	= 'h62;
		virtual_vram[ 17'h074CC ]	= 'h62;
		virtual_vram[ 17'h074CD ]	= 'h62;
		virtual_vram[ 17'h074CE ]	= 'h62;
		virtual_vram[ 17'h074CF ]	= 'h62;
		virtual_vram[ 17'h074D0 ]	= 'h62;
		virtual_vram[ 17'h074D1 ]	= 'h62;
		virtual_vram[ 17'h074D2 ]	= 'h62;
		virtual_vram[ 17'h074D3 ]	= 'h62;
		virtual_vram[ 17'h074D4 ]	= 'h62;
		virtual_vram[ 17'h074D5 ]	= 'h62;
		virtual_vram[ 17'h074D6 ]	= 'h62;
		virtual_vram[ 17'h074D7 ]	= 'h62;
		virtual_vram[ 17'h074D8 ]	= 'h62;
		virtual_vram[ 17'h074D9 ]	= 'h62;
		virtual_vram[ 17'h074DA ]	= 'h62;
		virtual_vram[ 17'h074DB ]	= 'h62;
		virtual_vram[ 17'h074DC ]	= 'h62;
		virtual_vram[ 17'h074DD ]	= 'h62;
		virtual_vram[ 17'h074DE ]	= 'h62;
		virtual_vram[ 17'h074DF ]	= 'h62;
		virtual_vram[ 17'h074E0 ]	= 'h62;
		virtual_vram[ 17'h074E1 ]	= 'h62;
		virtual_vram[ 17'h074E2 ]	= 'h62;
		virtual_vram[ 17'h074E3 ]	= 'h62;
		virtual_vram[ 17'h074E4 ]	= 'h62;
		virtual_vram[ 17'h074E5 ]	= 'h62;
		virtual_vram[ 17'h074E6 ]	= 'h62;
		virtual_vram[ 17'h074E7 ]	= 'h62;
		virtual_vram[ 17'h074E8 ]	= 'h62;
		virtual_vram[ 17'h074E9 ]	= 'h62;
		virtual_vram[ 17'h074EA ]	= 'h62;
		virtual_vram[ 17'h074EB ]	= 'h62;
		virtual_vram[ 17'h074EC ]	= 'h62;
		virtual_vram[ 17'h074ED ]	= 'h62;
		virtual_vram[ 17'h074EE ]	= 'h62;
		virtual_vram[ 17'h074EF ]	= 'h62;
		virtual_vram[ 17'h074F0 ]	= 'h62;
		virtual_vram[ 17'h074F1 ]	= 'h62;
		virtual_vram[ 17'h074F2 ]	= 'h62;
		virtual_vram[ 17'h074F3 ]	= 'h62;
		virtual_vram[ 17'h074F4 ]	= 'h62;
		virtual_vram[ 17'h074F5 ]	= 'h62;
		virtual_vram[ 17'h074F6 ]	= 'h62;
		virtual_vram[ 17'h074F7 ]	= 'h62;
		virtual_vram[ 17'h074F8 ]	= 'h62;
		virtual_vram[ 17'h074F9 ]	= 'h62;
		virtual_vram[ 17'h074FA ]	= 'h62;
		virtual_vram[ 17'h074FB ]	= 'h62;
		virtual_vram[ 17'h074FC ]	= 'h62;
		virtual_vram[ 17'h074FD ]	= 'h62;
		virtual_vram[ 17'h074FE ]	= 'h62;
		virtual_vram[ 17'h074FF ]	= 'h62;
		virtual_vram[ 17'h07500 ]	= 'h62;
		virtual_vram[ 17'h07501 ]	= 'h62;
		virtual_vram[ 17'h07502 ]	= 'h62;
		virtual_vram[ 17'h07503 ]	= 'h62;
		virtual_vram[ 17'h07504 ]	= 'h62;
		virtual_vram[ 17'h07505 ]	= 'h62;
		virtual_vram[ 17'h07506 ]	= 'h62;
		virtual_vram[ 17'h07507 ]	= 'h62;
		virtual_vram[ 17'h07508 ]	= 'h62;
		virtual_vram[ 17'h07509 ]	= 'h62;
		virtual_vram[ 17'h0750A ]	= 'h62;
		virtual_vram[ 17'h0750B ]	= 'h62;
		virtual_vram[ 17'h0750C ]	= 'h62;
		virtual_vram[ 17'h0750D ]	= 'h62;
		virtual_vram[ 17'h0750E ]	= 'h62;
		virtual_vram[ 17'h0750F ]	= 'h62;
		virtual_vram[ 17'h07510 ]	= 'h62;
		virtual_vram[ 17'h07511 ]	= 'h62;
		virtual_vram[ 17'h07512 ]	= 'h62;
		virtual_vram[ 17'h07513 ]	= 'h62;
		virtual_vram[ 17'h07514 ]	= 'h62;
		virtual_vram[ 17'h07515 ]	= 'h62;
		virtual_vram[ 17'h07516 ]	= 'h62;
		virtual_vram[ 17'h07517 ]	= 'h62;
		virtual_vram[ 17'h07518 ]	= 'h62;
		virtual_vram[ 17'h07519 ]	= 'h62;
		virtual_vram[ 17'h0751A ]	= 'h62;
		virtual_vram[ 17'h0751B ]	= 'h62;
		virtual_vram[ 17'h0751C ]	= 'h62;
		virtual_vram[ 17'h0751D ]	= 'h62;
		virtual_vram[ 17'h0751E ]	= 'h62;
		virtual_vram[ 17'h0751F ]	= 'h62;
		virtual_vram[ 17'h07520 ]	= 'h62;
		virtual_vram[ 17'h07521 ]	= 'h62;
		virtual_vram[ 17'h07522 ]	= 'h62;
		virtual_vram[ 17'h07523 ]	= 'h62;
		virtual_vram[ 17'h07524 ]	= 'h62;
		virtual_vram[ 17'h07525 ]	= 'h62;
		virtual_vram[ 17'h07526 ]	= 'h62;
		virtual_vram[ 17'h07527 ]	= 'h62;
		virtual_vram[ 17'h07528 ]	= 'h62;
		virtual_vram[ 17'h07529 ]	= 'h62;
		virtual_vram[ 17'h0752A ]	= 'h62;
		virtual_vram[ 17'h0752B ]	= 'h62;
		virtual_vram[ 17'h0752C ]	= 'h62;
		virtual_vram[ 17'h0752D ]	= 'h62;
		virtual_vram[ 17'h0752E ]	= 'h62;
		virtual_vram[ 17'h0752F ]	= 'h62;
		virtual_vram[ 17'h07530 ]	= 'h62;
		virtual_vram[ 17'h07531 ]	= 'h62;
		virtual_vram[ 17'h07532 ]	= 'h62;
		virtual_vram[ 17'h07533 ]	= 'h62;
		virtual_vram[ 17'h07534 ]	= 'h62;
		virtual_vram[ 17'h07535 ]	= 'h62;
		virtual_vram[ 17'h07536 ]	= 'h62;
		virtual_vram[ 17'h07537 ]	= 'h62;
		virtual_vram[ 17'h07538 ]	= 'h62;
		virtual_vram[ 17'h07539 ]	= 'h62;
		virtual_vram[ 17'h0753A ]	= 'h62;
		virtual_vram[ 17'h0753B ]	= 'h62;
		virtual_vram[ 17'h0753C ]	= 'h62;
		virtual_vram[ 17'h0753D ]	= 'h62;
		virtual_vram[ 17'h0753E ]	= 'h62;
		virtual_vram[ 17'h0753F ]	= 'h62;
		virtual_vram[ 17'h07540 ]	= 'h62;
		virtual_vram[ 17'h07541 ]	= 'h62;
		virtual_vram[ 17'h07542 ]	= 'h62;
		virtual_vram[ 17'h07543 ]	= 'h62;
		virtual_vram[ 17'h07544 ]	= 'h62;
		virtual_vram[ 17'h07545 ]	= 'h62;
		virtual_vram[ 17'h07546 ]	= 'h62;
		virtual_vram[ 17'h07547 ]	= 'h62;
		virtual_vram[ 17'h07548 ]	= 'h62;
		virtual_vram[ 17'h07549 ]	= 'h62;
		virtual_vram[ 17'h0754A ]	= 'h62;
		virtual_vram[ 17'h0754B ]	= 'h62;
		virtual_vram[ 17'h0754C ]	= 'h62;
		virtual_vram[ 17'h0754D ]	= 'h62;
		virtual_vram[ 17'h0754E ]	= 'h62;
		virtual_vram[ 17'h0754F ]	= 'h62;
		virtual_vram[ 17'h07550 ]	= 'h62;
		virtual_vram[ 17'h07551 ]	= 'h62;
		virtual_vram[ 17'h07552 ]	= 'h62;
		virtual_vram[ 17'h07553 ]	= 'h62;
		virtual_vram[ 17'h07554 ]	= 'h62;
		virtual_vram[ 17'h07555 ]	= 'h62;
		virtual_vram[ 17'h07556 ]	= 'h62;
		virtual_vram[ 17'h07557 ]	= 'h62;
		virtual_vram[ 17'h07558 ]	= 'h62;
		virtual_vram[ 17'h07559 ]	= 'h62;
		virtual_vram[ 17'h0755A ]	= 'h62;
		virtual_vram[ 17'h0755B ]	= 'h62;
		virtual_vram[ 17'h0755C ]	= 'h62;
		virtual_vram[ 17'h0755D ]	= 'h62;
		virtual_vram[ 17'h0755E ]	= 'h62;
		virtual_vram[ 17'h0755F ]	= 'h62;
		virtual_vram[ 17'h07560 ]	= 'h00;
		virtual_vram[ 17'h07561 ]	= 'h00;
		virtual_vram[ 17'h07562 ]	= 'h00;
		virtual_vram[ 17'h07563 ]	= 'h00;
		virtual_vram[ 17'h07564 ]	= 'h00;
		virtual_vram[ 17'h07565 ]	= 'h00;
		virtual_vram[ 17'h07566 ]	= 'h00;
		virtual_vram[ 17'h07567 ]	= 'h00;
		virtual_vram[ 17'h07568 ]	= 'h00;
		virtual_vram[ 17'h07569 ]	= 'h00;
		virtual_vram[ 17'h0756A ]	= 'h00;
		virtual_vram[ 17'h0756B ]	= 'h00;
		virtual_vram[ 17'h0756C ]	= 'h00;
		virtual_vram[ 17'h0756D ]	= 'h00;
		virtual_vram[ 17'h0756E ]	= 'h00;
		virtual_vram[ 17'h0756F ]	= 'h00;
		virtual_vram[ 17'h07570 ]	= 'h00;
		virtual_vram[ 17'h07571 ]	= 'h00;
		virtual_vram[ 17'h07572 ]	= 'h00;
		virtual_vram[ 17'h07573 ]	= 'h00;
		virtual_vram[ 17'h07574 ]	= 'h00;
		virtual_vram[ 17'h07575 ]	= 'h00;
		virtual_vram[ 17'h07576 ]	= 'h00;
		virtual_vram[ 17'h07577 ]	= 'h00;
		virtual_vram[ 17'h07578 ]	= 'h00;
		virtual_vram[ 17'h07579 ]	= 'h00;
		virtual_vram[ 17'h0757A ]	= 'h00;
		virtual_vram[ 17'h0757B ]	= 'h00;
		virtual_vram[ 17'h0757C ]	= 'h00;
		virtual_vram[ 17'h0757D ]	= 'h00;
		virtual_vram[ 17'h0757E ]	= 'h00;
		virtual_vram[ 17'h0757F ]	= 'h00;
		virtual_vram[ 17'h07580 ]	= 'h00;
		virtual_vram[ 17'h07581 ]	= 'h00;
		virtual_vram[ 17'h07582 ]	= 'h00;
		virtual_vram[ 17'h07583 ]	= 'h00;
		virtual_vram[ 17'h07584 ]	= 'h00;
		virtual_vram[ 17'h07585 ]	= 'h00;
		virtual_vram[ 17'h07586 ]	= 'h00;
		virtual_vram[ 17'h07587 ]	= 'h00;
		virtual_vram[ 17'h07588 ]	= 'h00;
		virtual_vram[ 17'h07589 ]	= 'h00;
		virtual_vram[ 17'h0758A ]	= 'h00;
		virtual_vram[ 17'h0758B ]	= 'h00;
		virtual_vram[ 17'h0758C ]	= 'h00;
		virtual_vram[ 17'h0758D ]	= 'h00;
		virtual_vram[ 17'h0758E ]	= 'h00;
		virtual_vram[ 17'h0758F ]	= 'h00;
		virtual_vram[ 17'h07590 ]	= 'h00;
		virtual_vram[ 17'h07591 ]	= 'h00;
		virtual_vram[ 17'h07592 ]	= 'h00;
		virtual_vram[ 17'h07593 ]	= 'h00;
		virtual_vram[ 17'h07594 ]	= 'h00;
		virtual_vram[ 17'h07595 ]	= 'h00;
		virtual_vram[ 17'h07596 ]	= 'h00;
		virtual_vram[ 17'h07597 ]	= 'h00;
		virtual_vram[ 17'h07598 ]	= 'h00;
		virtual_vram[ 17'h07599 ]	= 'h00;
		virtual_vram[ 17'h0759A ]	= 'h00;
		virtual_vram[ 17'h0759B ]	= 'h00;
		virtual_vram[ 17'h0759C ]	= 'h00;
		virtual_vram[ 17'h0759D ]	= 'h00;
		virtual_vram[ 17'h0759E ]	= 'h00;
		virtual_vram[ 17'h0759F ]	= 'h00;
		virtual_vram[ 17'h075A0 ]	= 'h00;
		virtual_vram[ 17'h075A1 ]	= 'h00;
		virtual_vram[ 17'h075A2 ]	= 'h00;
		virtual_vram[ 17'h075A3 ]	= 'h00;
		virtual_vram[ 17'h075A4 ]	= 'h00;
		virtual_vram[ 17'h075A5 ]	= 'h00;
		virtual_vram[ 17'h075A6 ]	= 'h00;
		virtual_vram[ 17'h075A7 ]	= 'h00;
		virtual_vram[ 17'h075A8 ]	= 'h00;
		virtual_vram[ 17'h075A9 ]	= 'h00;
		virtual_vram[ 17'h075AA ]	= 'h00;
		virtual_vram[ 17'h075AB ]	= 'h00;
		virtual_vram[ 17'h075AC ]	= 'h00;
		virtual_vram[ 17'h075AD ]	= 'h00;
		virtual_vram[ 17'h075AE ]	= 'h00;
		virtual_vram[ 17'h075AF ]	= 'h00;
		virtual_vram[ 17'h075B0 ]	= 'h00;
		virtual_vram[ 17'h075B1 ]	= 'h00;
		virtual_vram[ 17'h075B2 ]	= 'h00;
		virtual_vram[ 17'h075B3 ]	= 'h00;
		virtual_vram[ 17'h075B4 ]	= 'h00;
		virtual_vram[ 17'h075B5 ]	= 'h00;
		virtual_vram[ 17'h075B6 ]	= 'h00;
		virtual_vram[ 17'h075B7 ]	= 'h00;
		virtual_vram[ 17'h075B8 ]	= 'h00;
		virtual_vram[ 17'h075B9 ]	= 'h00;
		virtual_vram[ 17'h075BA ]	= 'h00;
		virtual_vram[ 17'h075BB ]	= 'h00;
		virtual_vram[ 17'h075BC ]	= 'h00;
		virtual_vram[ 17'h075BD ]	= 'h00;
		virtual_vram[ 17'h075BE ]	= 'h00;
		virtual_vram[ 17'h075BF ]	= 'h00;
		virtual_vram[ 17'h075C0 ]	= 'h00;
		virtual_vram[ 17'h075C1 ]	= 'h00;
		virtual_vram[ 17'h075C2 ]	= 'h00;
		virtual_vram[ 17'h075C3 ]	= 'h00;
		virtual_vram[ 17'h075C4 ]	= 'h00;
		virtual_vram[ 17'h075C5 ]	= 'h00;
		virtual_vram[ 17'h075C6 ]	= 'h00;
		virtual_vram[ 17'h075C7 ]	= 'h00;
		virtual_vram[ 17'h075C8 ]	= 'h00;
		virtual_vram[ 17'h075C9 ]	= 'h00;
		virtual_vram[ 17'h075CA ]	= 'h00;
		virtual_vram[ 17'h075CB ]	= 'h00;
		virtual_vram[ 17'h075CC ]	= 'h00;
		virtual_vram[ 17'h075CD ]	= 'h00;
		virtual_vram[ 17'h075CE ]	= 'h00;
		virtual_vram[ 17'h075CF ]	= 'h00;
		virtual_vram[ 17'h075D0 ]	= 'h00;
		virtual_vram[ 17'h075D1 ]	= 'h00;
		virtual_vram[ 17'h075D2 ]	= 'h00;
		virtual_vram[ 17'h075D3 ]	= 'h00;
		virtual_vram[ 17'h075D4 ]	= 'h00;
		virtual_vram[ 17'h075D5 ]	= 'h00;
		virtual_vram[ 17'h075D6 ]	= 'h00;
		virtual_vram[ 17'h075D7 ]	= 'h00;
		virtual_vram[ 17'h075D8 ]	= 'h00;
		virtual_vram[ 17'h075D9 ]	= 'h00;
		virtual_vram[ 17'h075DA ]	= 'h00;
		virtual_vram[ 17'h075DB ]	= 'h00;
		virtual_vram[ 17'h075DC ]	= 'h00;
		virtual_vram[ 17'h075DD ]	= 'h00;
		virtual_vram[ 17'h075DE ]	= 'h00;
		virtual_vram[ 17'h075DF ]	= 'h00;
		virtual_vram[ 17'h075E0 ]	= 'h00;
		virtual_vram[ 17'h075E1 ]	= 'h00;
		virtual_vram[ 17'h075E2 ]	= 'h00;
		virtual_vram[ 17'h075E3 ]	= 'h00;
		virtual_vram[ 17'h075E4 ]	= 'h00;
		virtual_vram[ 17'h075E5 ]	= 'h00;
		virtual_vram[ 17'h075E6 ]	= 'h00;
		virtual_vram[ 17'h075E7 ]	= 'h00;
		virtual_vram[ 17'h075E8 ]	= 'h00;
		virtual_vram[ 17'h075E9 ]	= 'h00;
		virtual_vram[ 17'h075EA ]	= 'h00;
		virtual_vram[ 17'h075EB ]	= 'h00;
		virtual_vram[ 17'h075EC ]	= 'h00;
		virtual_vram[ 17'h075ED ]	= 'h00;
		virtual_vram[ 17'h075EE ]	= 'h00;
		virtual_vram[ 17'h075EF ]	= 'h00;
		virtual_vram[ 17'h075F0 ]	= 'h00;
		virtual_vram[ 17'h075F1 ]	= 'h00;
		virtual_vram[ 17'h075F2 ]	= 'h00;
		virtual_vram[ 17'h075F3 ]	= 'h00;
		virtual_vram[ 17'h075F4 ]	= 'h00;
		virtual_vram[ 17'h075F5 ]	= 'h00;
		virtual_vram[ 17'h075F6 ]	= 'h00;
		virtual_vram[ 17'h075F7 ]	= 'h00;
		virtual_vram[ 17'h075F8 ]	= 'h00;
		virtual_vram[ 17'h075F9 ]	= 'h00;
		virtual_vram[ 17'h075FA ]	= 'h00;
		virtual_vram[ 17'h075FB ]	= 'h00;
		virtual_vram[ 17'h075FC ]	= 'h00;
		virtual_vram[ 17'h075FD ]	= 'h00;
		virtual_vram[ 17'h075FE ]	= 'h00;
		virtual_vram[ 17'h075FF ]	= 'h00;

		virtual_vram[ 17'h07600 ]	= 'h1F;
		virtual_vram[ 17'h07601 ]	= 'h58;
		virtual_vram[ 17'h07602 ]	= 'h00;
		virtual_vram[ 17'h07603 ]	= 'h00;
		virtual_vram[ 17'h07604 ]	= 'h1F;
		virtual_vram[ 17'h07605 ]	= 'h68;
		virtual_vram[ 17'h07606 ]	= 'h08;
		virtual_vram[ 17'h07607 ]	= 'h00;
		virtual_vram[ 17'h07608 ]	= 'h2F;
		virtual_vram[ 17'h07609 ]	= 'h58;
		virtual_vram[ 17'h0760A ]	= 'h10;
		virtual_vram[ 17'h0760B ]	= 'h00;
		virtual_vram[ 17'h0760C ]	= 'h2F;
		virtual_vram[ 17'h0760D ]	= 'h68;
		virtual_vram[ 17'h0760E ]	= 'h18;
		virtual_vram[ 17'h0760F ]	= 'h00;
		virtual_vram[ 17'h07610 ]	= 'h3F;
		virtual_vram[ 17'h07611 ]	= 'h58;
		virtual_vram[ 17'h07612 ]	= 'h20;
		virtual_vram[ 17'h07613 ]	= 'h00;
		virtual_vram[ 17'h07614 ]	= 'h3F;
		virtual_vram[ 17'h07615 ]	= 'h68;
		virtual_vram[ 17'h07616 ]	= 'h28;
		virtual_vram[ 17'h07617 ]	= 'h00;
		virtual_vram[ 17'h07618 ]	= 'h1F;
		virtual_vram[ 17'h07619 ]	= 'h78;
		virtual_vram[ 17'h0761A ]	= 'h30;
		virtual_vram[ 17'h0761B ]	= 'h00;
		virtual_vram[ 17'h0761C ]	= 'h1F;
		virtual_vram[ 17'h0761D ]	= 'h88;
		virtual_vram[ 17'h0761E ]	= 'h38;
		virtual_vram[ 17'h0761F ]	= 'h00;
		virtual_vram[ 17'h07620 ]	= 'h2F;
		virtual_vram[ 17'h07621 ]	= 'h78;
		virtual_vram[ 17'h07622 ]	= 'h40;
		virtual_vram[ 17'h07623 ]	= 'h00;
		virtual_vram[ 17'h07624 ]	= 'h2F;
		virtual_vram[ 17'h07625 ]	= 'h88;
		virtual_vram[ 17'h07626 ]	= 'h48;
		virtual_vram[ 17'h07627 ]	= 'h00;
		virtual_vram[ 17'h07628 ]	= 'h3F;
		virtual_vram[ 17'h07629 ]	= 'h88;
		virtual_vram[ 17'h0762A ]	= 'h50;
		virtual_vram[ 17'h0762B ]	= 'h00;
		virtual_vram[ 17'h0762C ]	= 'h1F;
		virtual_vram[ 17'h0762D ]	= 'h58;
		virtual_vram[ 17'h0762E ]	= 'h04;
		virtual_vram[ 17'h0762F ]	= 'h00;
		virtual_vram[ 17'h07630 ]	= 'h1F;
		virtual_vram[ 17'h07631 ]	= 'h68;
		virtual_vram[ 17'h07632 ]	= 'h0C;
		virtual_vram[ 17'h07633 ]	= 'h00;
		virtual_vram[ 17'h07634 ]	= 'h2F;
		virtual_vram[ 17'h07635 ]	= 'h58;
		virtual_vram[ 17'h07636 ]	= 'h14;
		virtual_vram[ 17'h07637 ]	= 'h00;
		virtual_vram[ 17'h07638 ]	= 'h2F;
		virtual_vram[ 17'h07639 ]	= 'h68;
		virtual_vram[ 17'h0763A ]	= 'h1C;
		virtual_vram[ 17'h0763B ]	= 'h00;
		virtual_vram[ 17'h0763C ]	= 'h3F;
		virtual_vram[ 17'h0763D ]	= 'h58;
		virtual_vram[ 17'h0763E ]	= 'h24;
		virtual_vram[ 17'h0763F ]	= 'h00;
		virtual_vram[ 17'h07640 ]	= 'h3F;
		virtual_vram[ 17'h07641 ]	= 'h68;
		virtual_vram[ 17'h07642 ]	= 'h2C;
		virtual_vram[ 17'h07643 ]	= 'h00;
		virtual_vram[ 17'h07644 ]	= 'h1F;
		virtual_vram[ 17'h07645 ]	= 'h78;
		virtual_vram[ 17'h07646 ]	= 'h34;
		virtual_vram[ 17'h07647 ]	= 'h00;
		virtual_vram[ 17'h07648 ]	= 'h1F;
		virtual_vram[ 17'h07649 ]	= 'h88;
		virtual_vram[ 17'h0764A ]	= 'h3C;
		virtual_vram[ 17'h0764B ]	= 'h00;
		virtual_vram[ 17'h0764C ]	= 'h2F;
		virtual_vram[ 17'h0764D ]	= 'h78;
		virtual_vram[ 17'h0764E ]	= 'h44;
		virtual_vram[ 17'h0764F ]	= 'h00;
		virtual_vram[ 17'h07650 ]	= 'h2F;
		virtual_vram[ 17'h07651 ]	= 'h88;
		virtual_vram[ 17'h07652 ]	= 'h4C;
		virtual_vram[ 17'h07653 ]	= 'h00;
		virtual_vram[ 17'h07654 ]	= 'hF5;
		virtual_vram[ 17'h07655 ]	= 'hC5;
		virtual_vram[ 17'h07656 ]	= 'hD5;
		virtual_vram[ 17'h07657 ]	= 'hE5;
		virtual_vram[ 17'h07658 ]	= 'hD8;
		virtual_vram[ 17'h07659 ]	= 'hD8;
		virtual_vram[ 17'h0765A ]	= 'hD8;
		virtual_vram[ 17'h0765B ]	= 'hD8;
		virtual_vram[ 17'h0765C ]	= 'hD8;
		virtual_vram[ 17'h0765D ]	= 'hD8;
		virtual_vram[ 17'h0765E ]	= 'hD8;
		virtual_vram[ 17'h0765F ]	= 'hD8;
		virtual_vram[ 17'h07660 ]	= 'hD8;
		virtual_vram[ 17'h07661 ]	= 'hD8;
		virtual_vram[ 17'h07662 ]	= 'hD8;
		virtual_vram[ 17'h07663 ]	= 'hD8;
		virtual_vram[ 17'h07664 ]	= 'hD8;
		virtual_vram[ 17'h07665 ]	= 'hD8;
		virtual_vram[ 17'h07666 ]	= 'hD8;
		virtual_vram[ 17'h07667 ]	= 'hD8;
		virtual_vram[ 17'h07668 ]	= 'hD8;
		virtual_vram[ 17'h07669 ]	= 'hD8;
		virtual_vram[ 17'h0766A ]	= 'hD8;
		virtual_vram[ 17'h0766B ]	= 'hD8;
		virtual_vram[ 17'h0766C ]	= 'hD8;
		virtual_vram[ 17'h0766D ]	= 'hD8;
		virtual_vram[ 17'h0766E ]	= 'hD8;
		virtual_vram[ 17'h0766F ]	= 'hD8;
		virtual_vram[ 17'h07670 ]	= 'hD8;
		virtual_vram[ 17'h07671 ]	= 'hD8;
		virtual_vram[ 17'h07672 ]	= 'hD8;
		virtual_vram[ 17'h07673 ]	= 'hD8;
		virtual_vram[ 17'h07674 ]	= 'hD8;
		virtual_vram[ 17'h07675 ]	= 'hD8;
		virtual_vram[ 17'h07676 ]	= 'hD8;
		virtual_vram[ 17'h07677 ]	= 'hD8;
		virtual_vram[ 17'h07678 ]	= 'hD8;
		virtual_vram[ 17'h07679 ]	= 'hD8;
		virtual_vram[ 17'h0767A ]	= 'hD8;
		virtual_vram[ 17'h0767B ]	= 'hD8;
		virtual_vram[ 17'h0767C ]	= 'hD8;
		virtual_vram[ 17'h0767D ]	= 'hD8;
		virtual_vram[ 17'h0767E ]	= 'hD8;
		virtual_vram[ 17'h0767F ]	= 'hD8;

		virtual_vram[ 17'h07800 ]	= 'h00;
		virtual_vram[ 17'h07801 ]	= 'h00;
		virtual_vram[ 17'h07802 ]	= 'h00;
		virtual_vram[ 17'h07803 ]	= 'h00;
		virtual_vram[ 17'h07804 ]	= 'h00;
		virtual_vram[ 17'h07805 ]	= 'h00;
		virtual_vram[ 17'h07806 ]	= 'h00;
		virtual_vram[ 17'h07807 ]	= 'h00;
		virtual_vram[ 17'h07808 ]	= 'hF0;
		virtual_vram[ 17'h07809 ]	= 'hFE;
		virtual_vram[ 17'h0780A ]	= 'hFE;
		virtual_vram[ 17'h0780B ]	= 'hFF;
		virtual_vram[ 17'h0780C ]	= 'hFF;
		virtual_vram[ 17'h0780D ]	= 'h77;
		virtual_vram[ 17'h0780E ]	= 'h77;
		virtual_vram[ 17'h0780F ]	= 'h73;
		virtual_vram[ 17'h07810 ]	= 'h00;
		virtual_vram[ 17'h07811 ]	= 'h00;
		virtual_vram[ 17'h07812 ]	= 'h00;
		virtual_vram[ 17'h07813 ]	= 'h00;
		virtual_vram[ 17'h07814 ]	= 'h00;
		virtual_vram[ 17'h07815 ]	= 'h00;
		virtual_vram[ 17'h07816 ]	= 'h00;
		virtual_vram[ 17'h07817 ]	= 'h00;
		virtual_vram[ 17'h07818 ]	= 'h00;
		virtual_vram[ 17'h07819 ]	= 'h00;
		virtual_vram[ 17'h0781A ]	= 'h03;
		virtual_vram[ 17'h0781B ]	= 'h07;
		virtual_vram[ 17'h0781C ]	= 'h0F;
		virtual_vram[ 17'h0781D ]	= 'h87;
		virtual_vram[ 17'h0781E ]	= 'h9B;
		virtual_vram[ 17'h0781F ]	= 'h8F;
		virtual_vram[ 17'h07820 ]	= 'h00;
		virtual_vram[ 17'h07821 ]	= 'h00;
		virtual_vram[ 17'h07822 ]	= 'h00;
		virtual_vram[ 17'h07823 ]	= 'h00;
		virtual_vram[ 17'h07824 ]	= 'h00;
		virtual_vram[ 17'h07825 ]	= 'h00;
		virtual_vram[ 17'h07826 ]	= 'h00;
		virtual_vram[ 17'h07827 ]	= 'h00;
		virtual_vram[ 17'h07828 ]	= 'h00;
		virtual_vram[ 17'h07829 ]	= 'h00;
		virtual_vram[ 17'h0782A ]	= 'h00;
		virtual_vram[ 17'h0782B ]	= 'h00;
		virtual_vram[ 17'h0782C ]	= 'h00;
		virtual_vram[ 17'h0782D ]	= 'h88;
		virtual_vram[ 17'h0782E ]	= 'h88;
		virtual_vram[ 17'h0782F ]	= 'h8C;
		virtual_vram[ 17'h07830 ]	= 'h00;
		virtual_vram[ 17'h07831 ]	= 'h00;
		virtual_vram[ 17'h07832 ]	= 'h00;
		virtual_vram[ 17'h07833 ]	= 'h00;
		virtual_vram[ 17'h07834 ]	= 'h00;
		virtual_vram[ 17'h07835 ]	= 'h00;
		virtual_vram[ 17'h07836 ]	= 'h00;
		virtual_vram[ 17'h07837 ]	= 'h00;
		virtual_vram[ 17'h07838 ]	= 'h00;
		virtual_vram[ 17'h07839 ]	= 'h00;
		virtual_vram[ 17'h0783A ]	= 'h00;
		virtual_vram[ 17'h0783B ]	= 'h00;
		virtual_vram[ 17'h0783C ]	= 'h00;
		virtual_vram[ 17'h0783D ]	= 'h78;
		virtual_vram[ 17'h0783E ]	= 'h64;
		virtual_vram[ 17'h0783F ]	= 'h70;
		virtual_vram[ 17'h07840 ]	= 'h00;
		virtual_vram[ 17'h07841 ]	= 'h00;
		virtual_vram[ 17'h07842 ]	= 'h00;
		virtual_vram[ 17'h07843 ]	= 'h00;
		virtual_vram[ 17'h07844 ]	= 'h00;
		virtual_vram[ 17'h07845 ]	= 'h00;
		virtual_vram[ 17'h07846 ]	= 'h00;
		virtual_vram[ 17'h07847 ]	= 'h00;
		virtual_vram[ 17'h07848 ]	= 'h00;
		virtual_vram[ 17'h07849 ]	= 'h00;
		virtual_vram[ 17'h0784A ]	= 'hF0;
		virtual_vram[ 17'h0784B ]	= 'hF8;
		virtual_vram[ 17'h0784C ]	= 'hF8;
		virtual_vram[ 17'h0784D ]	= 'hFC;
		virtual_vram[ 17'h0784E ]	= 'h3C;
		virtual_vram[ 17'h0784F ]	= 'h0E;
		virtual_vram[ 17'h07850 ]	= 'h00;
		virtual_vram[ 17'h07851 ]	= 'h00;
		virtual_vram[ 17'h07852 ]	= 'h00;
		virtual_vram[ 17'h07853 ]	= 'h00;
		virtual_vram[ 17'h07854 ]	= 'h00;
		virtual_vram[ 17'h07855 ]	= 'h00;
		virtual_vram[ 17'h07856 ]	= 'h00;
		virtual_vram[ 17'h07857 ]	= 'h00;
		virtual_vram[ 17'h07858 ]	= 'h00;
		virtual_vram[ 17'h07859 ]	= 'h00;
		virtual_vram[ 17'h0785A ]	= 'h00;
		virtual_vram[ 17'h0785B ]	= 'h7F;
		virtual_vram[ 17'h0785C ]	= 'h3F;
		virtual_vram[ 17'h0785D ]	= 'hBF;
		virtual_vram[ 17'h0785E ]	= 'hD3;
		virtual_vram[ 17'h0785F ]	= 'hF3;
		virtual_vram[ 17'h07860 ]	= 'h00;
		virtual_vram[ 17'h07861 ]	= 'h00;
		virtual_vram[ 17'h07862 ]	= 'h00;
		virtual_vram[ 17'h07863 ]	= 'h00;
		virtual_vram[ 17'h07864 ]	= 'h00;
		virtual_vram[ 17'h07865 ]	= 'h00;
		virtual_vram[ 17'h07866 ]	= 'h00;
		virtual_vram[ 17'h07867 ]	= 'h00;
		virtual_vram[ 17'h07868 ]	= 'h00;
		virtual_vram[ 17'h07869 ]	= 'h00;
		virtual_vram[ 17'h0786A ]	= 'h00;
		virtual_vram[ 17'h0786B ]	= 'h00;
		virtual_vram[ 17'h0786C ]	= 'h00;
		virtual_vram[ 17'h0786D ]	= 'h03;
		virtual_vram[ 17'h0786E ]	= 'hC3;
		virtual_vram[ 17'h0786F ]	= 'hF1;
		virtual_vram[ 17'h07870 ]	= 'h00;
		virtual_vram[ 17'h07871 ]	= 'h00;
		virtual_vram[ 17'h07872 ]	= 'h00;
		virtual_vram[ 17'h07873 ]	= 'h00;
		virtual_vram[ 17'h07874 ]	= 'h00;
		virtual_vram[ 17'h07875 ]	= 'h00;
		virtual_vram[ 17'h07876 ]	= 'h00;
		virtual_vram[ 17'h07877 ]	= 'h00;
		virtual_vram[ 17'h07878 ]	= 'h00;
		virtual_vram[ 17'h07879 ]	= 'h00;
		virtual_vram[ 17'h0787A ]	= 'h00;
		virtual_vram[ 17'h0787B ]	= 'h00;
		virtual_vram[ 17'h0787C ]	= 'hC0;
		virtual_vram[ 17'h0787D ]	= 'h40;
		virtual_vram[ 17'h0787E ]	= 'h2C;
		virtual_vram[ 17'h0787F ]	= 'h0C;
		virtual_vram[ 17'h07880 ]	= 'h73;
		virtual_vram[ 17'h07881 ]	= 'h7B;
		virtual_vram[ 17'h07882 ]	= 'h79;
		virtual_vram[ 17'h07883 ]	= 'h39;
		virtual_vram[ 17'h07884 ]	= 'h39;
		virtual_vram[ 17'h07885 ]	= 'h3C;
		virtual_vram[ 17'h07886 ]	= 'h3C;
		virtual_vram[ 17'h07887 ]	= 'h3C;
		virtual_vram[ 17'h07888 ]	= 'h3F;
		virtual_vram[ 17'h07889 ]	= 'h1B;
		virtual_vram[ 17'h0788A ]	= 'h1D;
		virtual_vram[ 17'h0788B ]	= 'h9D;
		virtual_vram[ 17'h0788C ]	= 'h9E;
		virtual_vram[ 17'h0788D ]	= 'h9F;
		virtual_vram[ 17'h0788E ]	= 'hCF;
		virtual_vram[ 17'h0788F ]	= 'hCF;
		virtual_vram[ 17'h07890 ]	= 'hCF;
		virtual_vram[ 17'h07891 ]	= 'h8F;
		virtual_vram[ 17'h07892 ]	= 'hC7;
		virtual_vram[ 17'h07893 ]	= 'hE7;
		virtual_vram[ 17'h07894 ]	= 'hE7;
		virtual_vram[ 17'h07895 ]	= 'hE7;
		virtual_vram[ 17'h07896 ]	= 'hF7;
		virtual_vram[ 17'h07897 ]	= 'hF3;
		virtual_vram[ 17'h07898 ]	= 'hF3;
		virtual_vram[ 17'h07899 ]	= 'hFB;
		virtual_vram[ 17'h0789A ]	= 'hFB;
		virtual_vram[ 17'h0789B ]	= 'hFB;
		virtual_vram[ 17'h0789C ]	= 'h3D;
		virtual_vram[ 17'h0789D ]	= 'h3C;
		virtual_vram[ 17'h0789E ]	= 'h1C;
		virtual_vram[ 17'h0789F ]	= 'h00;
		virtual_vram[ 17'h078A0 ]	= 'h8C;
		virtual_vram[ 17'h078A1 ]	= 'h84;
		virtual_vram[ 17'h078A2 ]	= 'h86;
		virtual_vram[ 17'h078A3 ]	= 'hC6;
		virtual_vram[ 17'h078A4 ]	= 'hC6;
		virtual_vram[ 17'h078A5 ]	= 'hC3;
		virtual_vram[ 17'h078A6 ]	= 'hC3;
		virtual_vram[ 17'h078A7 ]	= 'hC3;
		virtual_vram[ 17'h078A8 ]	= 'hC0;
		virtual_vram[ 17'h078A9 ]	= 'hE4;
		virtual_vram[ 17'h078AA ]	= 'hE2;
		virtual_vram[ 17'h078AB ]	= 'h62;
		virtual_vram[ 17'h078AC ]	= 'h61;
		virtual_vram[ 17'h078AD ]	= 'h60;
		virtual_vram[ 17'h078AE ]	= 'h30;
		virtual_vram[ 17'h078AF ]	= 'h30;
		virtual_vram[ 17'h078B0 ]	= 'h30;
		virtual_vram[ 17'h078B1 ]	= 'h70;
		virtual_vram[ 17'h078B2 ]	= 'h38;
		virtual_vram[ 17'h078B3 ]	= 'h18;
		virtual_vram[ 17'h078B4 ]	= 'h18;
		virtual_vram[ 17'h078B5 ]	= 'h18;
		virtual_vram[ 17'h078B6 ]	= 'h08;
		virtual_vram[ 17'h078B7 ]	= 'h0C;
		virtual_vram[ 17'h078B8 ]	= 'h0C;
		virtual_vram[ 17'h078B9 ]	= 'h04;
		virtual_vram[ 17'h078BA ]	= 'h04;
		virtual_vram[ 17'h078BB ]	= 'h04;
		virtual_vram[ 17'h078BC ]	= 'hC2;
		virtual_vram[ 17'h078BD ]	= 'hC3;
		virtual_vram[ 17'h078BE ]	= 'hE3;
		virtual_vram[ 17'h078BF ]	= 'hBF;
		virtual_vram[ 17'h078C0 ]	= 'h1E;
		virtual_vram[ 17'h078C1 ]	= 'h1E;
		virtual_vram[ 17'h078C2 ]	= 'h00;
		virtual_vram[ 17'h078C3 ]	= 'h00;
		virtual_vram[ 17'h078C4 ]	= 'hBE;
		virtual_vram[ 17'h078C5 ]	= 'hBE;
		virtual_vram[ 17'h078C6 ]	= 'hB6;
		virtual_vram[ 17'h078C7 ]	= 'h8F;
		virtual_vram[ 17'h078C8 ]	= 'hCF;
		virtual_vram[ 17'h078C9 ]	= 'hC7;
		virtual_vram[ 17'h078CA ]	= 'hE7;
		virtual_vram[ 17'h078CB ]	= 'hFF;
		virtual_vram[ 17'h078CC ]	= 'hEF;
		virtual_vram[ 17'h078CD ]	= 'h9E;
		virtual_vram[ 17'h078CE ]	= 'h7E;
		virtual_vram[ 17'h078CF ]	= 'h00;
		virtual_vram[ 17'h078D0 ]	= 'hF3;
		virtual_vram[ 17'h078D1 ]	= 'hF3;
		virtual_vram[ 17'h078D2 ]	= 'hF3;
		virtual_vram[ 17'h078D3 ]	= 'hF3;
		virtual_vram[ 17'h078D4 ]	= 'hF1;
		virtual_vram[ 17'h078D5 ]	= 'h79;
		virtual_vram[ 17'h078D6 ]	= 'h79;
		virtual_vram[ 17'h078D7 ]	= 'h79;
		virtual_vram[ 17'h078D8 ]	= 'h79;
		virtual_vram[ 17'h078D9 ]	= 'h79;
		virtual_vram[ 17'h078DA ]	= 'h79;
		virtual_vram[ 17'h078DB ]	= 'h5F;
		virtual_vram[ 17'h078DC ]	= 'h7F;
		virtual_vram[ 17'h078DD ]	= 'h1F;
		virtual_vram[ 17'h078DE ]	= 'h80;
		virtual_vram[ 17'h078DF ]	= 'h00;
		virtual_vram[ 17'h078E0 ]	= 'hE1;
		virtual_vram[ 17'h078E1 ]	= 'hE1;
		virtual_vram[ 17'h078E2 ]	= 'hDD;
		virtual_vram[ 17'h078E3 ]	= 'h3B;
		virtual_vram[ 17'h078E4 ]	= 'h41;
		virtual_vram[ 17'h078E5 ]	= 'h41;
		virtual_vram[ 17'h078E6 ]	= 'h49;
		virtual_vram[ 17'h078E7 ]	= 'h70;
		virtual_vram[ 17'h078E8 ]	= 'h30;
		virtual_vram[ 17'h078E9 ]	= 'h38;
		virtual_vram[ 17'h078EA ]	= 'h18;
		virtual_vram[ 17'h078EB ]	= 'h00;
		virtual_vram[ 17'h078EC ]	= 'h10;
		virtual_vram[ 17'h078ED ]	= 'h61;
		virtual_vram[ 17'h078EE ]	= 'h00;
		virtual_vram[ 17'h078EF ]	= 'hFC;
		virtual_vram[ 17'h078F0 ]	= 'h0C;
		virtual_vram[ 17'h078F1 ]	= 'h0C;
		virtual_vram[ 17'h078F2 ]	= 'h0C;
		virtual_vram[ 17'h078F3 ]	= 'h0C;
		virtual_vram[ 17'h078F4 ]	= 'h0E;
		virtual_vram[ 17'h078F5 ]	= 'h86;
		virtual_vram[ 17'h078F6 ]	= 'h86;
		virtual_vram[ 17'h078F7 ]	= 'h86;
		virtual_vram[ 17'h078F8 ]	= 'h86;
		virtual_vram[ 17'h078F9 ]	= 'h86;
		virtual_vram[ 17'h078FA ]	= 'h86;
		virtual_vram[ 17'h078FB ]	= 'hA0;
		virtual_vram[ 17'h078FC ]	= 'h80;
		virtual_vram[ 17'h078FD ]	= 'hE0;
		virtual_vram[ 17'h078FE ]	= 'h7F;
		virtual_vram[ 17'h078FF ]	= 'h7F;
		virtual_vram[ 17'h07900 ]	= 'hE0;
		virtual_vram[ 17'h07901 ]	= 'h00;
		virtual_vram[ 17'h07902 ]	= 'h00;
		virtual_vram[ 17'h07903 ]	= 'h00;
		virtual_vram[ 17'h07904 ]	= 'h00;
		virtual_vram[ 17'h07905 ]	= 'h00;
		virtual_vram[ 17'h07906 ]	= 'h00;
		virtual_vram[ 17'h07907 ]	= 'h00;
		virtual_vram[ 17'h07908 ]	= 'h00;
		virtual_vram[ 17'h07909 ]	= 'h00;
		virtual_vram[ 17'h0790A ]	= 'h00;
		virtual_vram[ 17'h0790B ]	= 'h00;
		virtual_vram[ 17'h0790C ]	= 'h00;
		virtual_vram[ 17'h0790D ]	= 'h00;
		virtual_vram[ 17'h0790E ]	= 'h00;
		virtual_vram[ 17'h0790F ]	= 'h00;
		virtual_vram[ 17'h07910 ]	= 'h00;
		virtual_vram[ 17'h07911 ]	= 'h00;
		virtual_vram[ 17'h07912 ]	= 'h00;
		virtual_vram[ 17'h07913 ]	= 'h00;
		virtual_vram[ 17'h07914 ]	= 'h00;
		virtual_vram[ 17'h07915 ]	= 'h00;
		virtual_vram[ 17'h07916 ]	= 'h00;
		virtual_vram[ 17'h07917 ]	= 'h00;
		virtual_vram[ 17'h07918 ]	= 'h00;
		virtual_vram[ 17'h07919 ]	= 'h00;
		virtual_vram[ 17'h0791A ]	= 'h00;
		virtual_vram[ 17'h0791B ]	= 'h00;
		virtual_vram[ 17'h0791C ]	= 'h00;
		virtual_vram[ 17'h0791D ]	= 'h00;
		virtual_vram[ 17'h0791E ]	= 'h00;
		virtual_vram[ 17'h0791F ]	= 'h00;
		virtual_vram[ 17'h07920 ]	= 'h1F;
		virtual_vram[ 17'h07921 ]	= 'hFC;
		virtual_vram[ 17'h07922 ]	= 'hFC;
		virtual_vram[ 17'h07923 ]	= 'h80;
		virtual_vram[ 17'h07924 ]	= 'h00;
		virtual_vram[ 17'h07925 ]	= 'h00;
		virtual_vram[ 17'h07926 ]	= 'h00;
		virtual_vram[ 17'h07927 ]	= 'h00;
		virtual_vram[ 17'h07928 ]	= 'h00;
		virtual_vram[ 17'h07929 ]	= 'h00;
		virtual_vram[ 17'h0792A ]	= 'h00;
		virtual_vram[ 17'h0792B ]	= 'h00;
		virtual_vram[ 17'h0792C ]	= 'h00;
		virtual_vram[ 17'h0792D ]	= 'h00;
		virtual_vram[ 17'h0792E ]	= 'h00;
		virtual_vram[ 17'h0792F ]	= 'h00;
		virtual_vram[ 17'h07930 ]	= 'h79;
		virtual_vram[ 17'h07931 ]	= 'hF0;
		virtual_vram[ 17'h07932 ]	= 'h00;
		virtual_vram[ 17'h07933 ]	= 'h00;
		virtual_vram[ 17'h07934 ]	= 'h00;
		virtual_vram[ 17'h07935 ]	= 'h00;
		virtual_vram[ 17'h07936 ]	= 'h00;
		virtual_vram[ 17'h07937 ]	= 'h00;
		virtual_vram[ 17'h07938 ]	= 'h00;
		virtual_vram[ 17'h07939 ]	= 'h00;
		virtual_vram[ 17'h0793A ]	= 'h00;
		virtual_vram[ 17'h0793B ]	= 'h00;
		virtual_vram[ 17'h0793C ]	= 'h00;
		virtual_vram[ 17'h0793D ]	= 'h00;
		virtual_vram[ 17'h0793E ]	= 'h00;
		virtual_vram[ 17'h0793F ]	= 'h00;
		virtual_vram[ 17'h07940 ]	= 'h00;
		virtual_vram[ 17'h07941 ]	= 'h00;
		virtual_vram[ 17'h07942 ]	= 'h00;
		virtual_vram[ 17'h07943 ]	= 'h00;
		virtual_vram[ 17'h07944 ]	= 'h00;
		virtual_vram[ 17'h07945 ]	= 'h00;
		virtual_vram[ 17'h07946 ]	= 'h00;
		virtual_vram[ 17'h07947 ]	= 'h00;
		virtual_vram[ 17'h07948 ]	= 'h00;
		virtual_vram[ 17'h07949 ]	= 'h00;
		virtual_vram[ 17'h0794A ]	= 'h00;
		virtual_vram[ 17'h0794B ]	= 'h00;
		virtual_vram[ 17'h0794C ]	= 'h00;
		virtual_vram[ 17'h0794D ]	= 'h00;
		virtual_vram[ 17'h0794E ]	= 'h00;
		virtual_vram[ 17'h0794F ]	= 'h00;
		virtual_vram[ 17'h07950 ]	= 'h00;
		virtual_vram[ 17'h07951 ]	= 'h00;
		virtual_vram[ 17'h07952 ]	= 'h00;
		virtual_vram[ 17'h07953 ]	= 'h00;
		virtual_vram[ 17'h07954 ]	= 'h00;
		virtual_vram[ 17'h07955 ]	= 'h00;
		virtual_vram[ 17'h07956 ]	= 'h00;
		virtual_vram[ 17'h07957 ]	= 'h00;
		virtual_vram[ 17'h07958 ]	= 'h00;
		virtual_vram[ 17'h07959 ]	= 'h00;
		virtual_vram[ 17'h0795A ]	= 'h00;
		virtual_vram[ 17'h0795B ]	= 'h00;
		virtual_vram[ 17'h0795C ]	= 'h00;
		virtual_vram[ 17'h0795D ]	= 'h00;
		virtual_vram[ 17'h0795E ]	= 'h00;
		virtual_vram[ 17'h0795F ]	= 'h00;
		virtual_vram[ 17'h07960 ]	= 'hFE;
		virtual_vram[ 17'h07961 ]	= 'h00;
		virtual_vram[ 17'h07962 ]	= 'h00;
		virtual_vram[ 17'h07963 ]	= 'h00;
		virtual_vram[ 17'h07964 ]	= 'h00;
		virtual_vram[ 17'h07965 ]	= 'h00;
		virtual_vram[ 17'h07966 ]	= 'h00;
		virtual_vram[ 17'h07967 ]	= 'h00;
		virtual_vram[ 17'h07968 ]	= 'h00;
		virtual_vram[ 17'h07969 ]	= 'h00;
		virtual_vram[ 17'h0796A ]	= 'h00;
		virtual_vram[ 17'h0796B ]	= 'h00;
		virtual_vram[ 17'h0796C ]	= 'h00;
		virtual_vram[ 17'h0796D ]	= 'h00;
		virtual_vram[ 17'h0796E ]	= 'h00;
		virtual_vram[ 17'h0796F ]	= 'h00;
		virtual_vram[ 17'h07970 ]	= 'h00;
		virtual_vram[ 17'h07971 ]	= 'h00;
		virtual_vram[ 17'h07972 ]	= 'h00;
		virtual_vram[ 17'h07973 ]	= 'h00;
		virtual_vram[ 17'h07974 ]	= 'h00;
		virtual_vram[ 17'h07975 ]	= 'h00;
		virtual_vram[ 17'h07976 ]	= 'h00;
		virtual_vram[ 17'h07977 ]	= 'h00;
		virtual_vram[ 17'h07978 ]	= 'h00;
		virtual_vram[ 17'h07979 ]	= 'h00;
		virtual_vram[ 17'h0797A ]	= 'h00;
		virtual_vram[ 17'h0797B ]	= 'h00;
		virtual_vram[ 17'h0797C ]	= 'h00;
		virtual_vram[ 17'h0797D ]	= 'h00;
		virtual_vram[ 17'h0797E ]	= 'h00;
		virtual_vram[ 17'h0797F ]	= 'h00;
		virtual_vram[ 17'h07980 ]	= 'h00;
		virtual_vram[ 17'h07981 ]	= 'h00;
		virtual_vram[ 17'h07982 ]	= 'h00;
		virtual_vram[ 17'h07983 ]	= 'h00;
		virtual_vram[ 17'h07984 ]	= 'h00;
		virtual_vram[ 17'h07985 ]	= 'h00;
		virtual_vram[ 17'h07986 ]	= 'h00;
		virtual_vram[ 17'h07987 ]	= 'h00;
		virtual_vram[ 17'h07988 ]	= 'h00;
		virtual_vram[ 17'h07989 ]	= 'h00;
		virtual_vram[ 17'h0798A ]	= 'h00;
		virtual_vram[ 17'h0798B ]	= 'h0C;
		virtual_vram[ 17'h0798C ]	= 'h1C;
		virtual_vram[ 17'h0798D ]	= 'h0C;
		virtual_vram[ 17'h0798E ]	= 'h96;
		virtual_vram[ 17'h0798F ]	= 'hDE;
		virtual_vram[ 17'h07990 ]	= 'h00;
		virtual_vram[ 17'h07991 ]	= 'h00;
		virtual_vram[ 17'h07992 ]	= 'h00;
		virtual_vram[ 17'h07993 ]	= 'h00;
		virtual_vram[ 17'h07994 ]	= 'h00;
		virtual_vram[ 17'h07995 ]	= 'h00;
		virtual_vram[ 17'h07996 ]	= 'h00;
		virtual_vram[ 17'h07997 ]	= 'h00;
		virtual_vram[ 17'h07998 ]	= 'h00;
		virtual_vram[ 17'h07999 ]	= 'h00;
		virtual_vram[ 17'h0799A ]	= 'h00;
		virtual_vram[ 17'h0799B ]	= 'hF8;
		virtual_vram[ 17'h0799C ]	= 'hF8;
		virtual_vram[ 17'h0799D ]	= 'hF8;
		virtual_vram[ 17'h0799E ]	= 'hF8;
		virtual_vram[ 17'h0799F ]	= 'hF8;
		virtual_vram[ 17'h079A0 ]	= 'h00;
		virtual_vram[ 17'h079A1 ]	= 'h00;
		virtual_vram[ 17'h079A2 ]	= 'h00;
		virtual_vram[ 17'h079A3 ]	= 'h00;
		virtual_vram[ 17'h079A4 ]	= 'h00;
		virtual_vram[ 17'h079A5 ]	= 'h00;
		virtual_vram[ 17'h079A6 ]	= 'h00;
		virtual_vram[ 17'h079A7 ]	= 'h00;
		virtual_vram[ 17'h079A8 ]	= 'h00;
		virtual_vram[ 17'h079A9 ]	= 'h00;
		virtual_vram[ 17'h079AA ]	= 'h00;
		virtual_vram[ 17'h079AB ]	= 'h00;
		virtual_vram[ 17'h079AC ]	= 'h00;
		virtual_vram[ 17'h079AD ]	= 'h00;
		virtual_vram[ 17'h079AE ]	= 'h00;
		virtual_vram[ 17'h079AF ]	= 'h00;
		virtual_vram[ 17'h079B0 ]	= 'h00;
		virtual_vram[ 17'h079B1 ]	= 'h00;
		virtual_vram[ 17'h079B2 ]	= 'h00;
		virtual_vram[ 17'h079B3 ]	= 'h00;
		virtual_vram[ 17'h079B4 ]	= 'h00;
		virtual_vram[ 17'h079B5 ]	= 'h00;
		virtual_vram[ 17'h079B6 ]	= 'h00;
		virtual_vram[ 17'h079B7 ]	= 'h00;
		virtual_vram[ 17'h079B8 ]	= 'h00;
		virtual_vram[ 17'h079B9 ]	= 'h00;
		virtual_vram[ 17'h079BA ]	= 'h00;
		virtual_vram[ 17'h079BB ]	= 'h00;
		virtual_vram[ 17'h079BC ]	= 'h00;
		virtual_vram[ 17'h079BD ]	= 'h00;
		virtual_vram[ 17'h079BE ]	= 'h00;
		virtual_vram[ 17'h079BF ]	= 'h00;
		virtual_vram[ 17'h079C0 ]	= 'h00;
		virtual_vram[ 17'h079C1 ]	= 'h00;
		virtual_vram[ 17'h079C2 ]	= 'h00;
		virtual_vram[ 17'h079C3 ]	= 'h00;
		virtual_vram[ 17'h079C4 ]	= 'h00;
		virtual_vram[ 17'h079C5 ]	= 'h00;
		virtual_vram[ 17'h079C6 ]	= 'h00;
		virtual_vram[ 17'h079C7 ]	= 'h00;
		virtual_vram[ 17'h079C8 ]	= 'h00;
		virtual_vram[ 17'h079C9 ]	= 'h00;
		virtual_vram[ 17'h079CA ]	= 'h3F;
		virtual_vram[ 17'h079CB ]	= 'h7F;
		virtual_vram[ 17'h079CC ]	= 'hBF;
		virtual_vram[ 17'h079CD ]	= 'hFE;
		virtual_vram[ 17'h079CE ]	= 'hF3;
		virtual_vram[ 17'h079CF ]	= 'hF3;
		virtual_vram[ 17'h079D0 ]	= 'h00;
		virtual_vram[ 17'h079D1 ]	= 'h00;
		virtual_vram[ 17'h079D2 ]	= 'h00;
		virtual_vram[ 17'h079D3 ]	= 'h00;
		virtual_vram[ 17'h079D4 ]	= 'h00;
		virtual_vram[ 17'h079D5 ]	= 'h00;
		virtual_vram[ 17'h079D6 ]	= 'h00;
		virtual_vram[ 17'h079D7 ]	= 'h00;
		virtual_vram[ 17'h079D8 ]	= 'h00;
		virtual_vram[ 17'h079D9 ]	= 'h00;
		virtual_vram[ 17'h079DA ]	= 'h07;
		virtual_vram[ 17'h079DB ]	= 'h8B;
		virtual_vram[ 17'h079DC ]	= 'h4F;
		virtual_vram[ 17'h079DD ]	= 'hCF;
		virtual_vram[ 17'h079DE ]	= 'h9E;
		virtual_vram[ 17'h079DF ]	= 'hDE;
		virtual_vram[ 17'h079E0 ]	= 'h00;
		virtual_vram[ 17'h079E1 ]	= 'h00;
		virtual_vram[ 17'h079E2 ]	= 'h00;
		virtual_vram[ 17'h079E3 ]	= 'h00;
		virtual_vram[ 17'h079E4 ]	= 'h00;
		virtual_vram[ 17'h079E5 ]	= 'h00;
		virtual_vram[ 17'h079E6 ]	= 'h00;
		virtual_vram[ 17'h079E7 ]	= 'h00;
		virtual_vram[ 17'h079E8 ]	= 'h00;
		virtual_vram[ 17'h079E9 ]	= 'h00;
		virtual_vram[ 17'h079EA ]	= 'h00;
		virtual_vram[ 17'h079EB ]	= 'h00;
		virtual_vram[ 17'h079EC ]	= 'h40;
		virtual_vram[ 17'h079ED ]	= 'h01;
		virtual_vram[ 17'h079EE ]	= 'h0C;
		virtual_vram[ 17'h079EF ]	= 'h0C;
		virtual_vram[ 17'h079F0 ]	= 'h00;
		virtual_vram[ 17'h079F1 ]	= 'h00;
		virtual_vram[ 17'h079F2 ]	= 'h00;
		virtual_vram[ 17'h079F3 ]	= 'h00;
		virtual_vram[ 17'h079F4 ]	= 'h00;
		virtual_vram[ 17'h079F5 ]	= 'h00;
		virtual_vram[ 17'h079F6 ]	= 'h00;
		virtual_vram[ 17'h079F7 ]	= 'h00;
		virtual_vram[ 17'h079F8 ]	= 'h00;
		virtual_vram[ 17'h079F9 ]	= 'h00;
		virtual_vram[ 17'h079FA ]	= 'h00;
		virtual_vram[ 17'h079FB ]	= 'h04;
		virtual_vram[ 17'h079FC ]	= 'hB0;
		virtual_vram[ 17'h079FD ]	= 'h30;
		virtual_vram[ 17'h079FE ]	= 'h61;
		virtual_vram[ 17'h079FF ]	= 'h21;
		virtual_vram[ 17'h07A00 ]	= 'hDE;
		virtual_vram[ 17'h07A01 ]	= 'h9F;
		virtual_vram[ 17'h07A02 ]	= 'h5F;
		virtual_vram[ 17'h07A03 ]	= 'hDF;
		virtual_vram[ 17'h07A04 ]	= 'hDF;
		virtual_vram[ 17'h07A05 ]	= 'hDF;
		virtual_vram[ 17'h07A06 ]	= 'hDF;
		virtual_vram[ 17'h07A07 ]	= 'hDF;
		virtual_vram[ 17'h07A08 ]	= 'hDD;
		virtual_vram[ 17'h07A09 ]	= 'hDC;
		virtual_vram[ 17'h07A0A ]	= 'hDC;
		virtual_vram[ 17'h07A0B ]	= 'hDC;
		virtual_vram[ 17'h07A0C ]	= 'hDC;
		virtual_vram[ 17'h07A0D ]	= 'h98;
		virtual_vram[ 17'h07A0E ]	= 'h00;
		virtual_vram[ 17'h07A0F ]	= 'h00;
		virtual_vram[ 17'h07A10 ]	= 'h79;
		virtual_vram[ 17'h07A11 ]	= 'h79;
		virtual_vram[ 17'h07A12 ]	= 'h79;
		virtual_vram[ 17'h07A13 ]	= 'h79;
		virtual_vram[ 17'h07A14 ]	= 'h39;
		virtual_vram[ 17'h07A15 ]	= 'hB9;
		virtual_vram[ 17'h07A16 ]	= 'hB9;
		virtual_vram[ 17'h07A17 ]	= 'hDB;
		virtual_vram[ 17'h07A18 ]	= 'hFB;
		virtual_vram[ 17'h07A19 ]	= 'hFB;
		virtual_vram[ 17'h07A1A ]	= 'hFB;
		virtual_vram[ 17'h07A1B ]	= 'hFB;
		virtual_vram[ 17'h07A1C ]	= 'h7A;
		virtual_vram[ 17'h07A1D ]	= 'h79;
		virtual_vram[ 17'h07A1E ]	= 'h00;
		virtual_vram[ 17'h07A1F ]	= 'h00;
		virtual_vram[ 17'h07A20 ]	= 'h21;
		virtual_vram[ 17'h07A21 ]	= 'h60;
		virtual_vram[ 17'h07A22 ]	= 'hA0;
		virtual_vram[ 17'h07A23 ]	= 'h20;
		virtual_vram[ 17'h07A24 ]	= 'h20;
		virtual_vram[ 17'h07A25 ]	= 'h20;
		virtual_vram[ 17'h07A26 ]	= 'h20;
		virtual_vram[ 17'h07A27 ]	= 'h20;
		virtual_vram[ 17'h07A28 ]	= 'h22;
		virtual_vram[ 17'h07A29 ]	= 'h23;
		virtual_vram[ 17'h07A2A ]	= 'h23;
		virtual_vram[ 17'h07A2B ]	= 'h23;
		virtual_vram[ 17'h07A2C ]	= 'h23;
		virtual_vram[ 17'h07A2D ]	= 'h67;
		virtual_vram[ 17'h07A2E ]	= 'h9E;
		virtual_vram[ 17'h07A2F ]	= 'h1E;
		virtual_vram[ 17'h07A30 ]	= 'h86;
		virtual_vram[ 17'h07A31 ]	= 'h86;
		virtual_vram[ 17'h07A32 ]	= 'h86;
		virtual_vram[ 17'h07A33 ]	= 'h86;
		virtual_vram[ 17'h07A34 ]	= 'hC6;
		virtual_vram[ 17'h07A35 ]	= 'h46;
		virtual_vram[ 17'h07A36 ]	= 'h46;
		virtual_vram[ 17'h07A37 ]	= 'h24;
		virtual_vram[ 17'h07A38 ]	= 'h04;
		virtual_vram[ 17'h07A39 ]	= 'h04;
		virtual_vram[ 17'h07A3A ]	= 'h04;
		virtual_vram[ 17'h07A3B ]	= 'h04;
		virtual_vram[ 17'h07A3C ]	= 'h85;
		virtual_vram[ 17'h07A3D ]	= 'h86;
		virtual_vram[ 17'h07A3E ]	= 'h7D;
		virtual_vram[ 17'h07A3F ]	= 'h78;
		virtual_vram[ 17'h07A40 ]	= 'hD3;
		virtual_vram[ 17'h07A41 ]	= 'hE3;
		virtual_vram[ 17'h07A42 ]	= 'hE7;
		virtual_vram[ 17'h07A43 ]	= 'hE7;
		virtual_vram[ 17'h07A44 ]	= 'hE7;
		virtual_vram[ 17'h07A45 ]	= 'hE7;
		virtual_vram[ 17'h07A46 ]	= 'hE7;
		virtual_vram[ 17'h07A47 ]	= 'hE7;
		virtual_vram[ 17'h07A48 ]	= 'hCF;
		virtual_vram[ 17'h07A49 ]	= 'hCF;
		virtual_vram[ 17'h07A4A ]	= 'hCF;
		virtual_vram[ 17'h07A4B ]	= 'hFE;
		virtual_vram[ 17'h07A4C ]	= 'hFE;
		virtual_vram[ 17'h07A4D ]	= 'hEC;
		virtual_vram[ 17'h07A4E ]	= 'hF0;
		virtual_vram[ 17'h07A4F ]	= 'hE0;
		virtual_vram[ 17'h07A50 ]	= 'hDE;
		virtual_vram[ 17'h07A51 ]	= 'hDE;
		virtual_vram[ 17'h07A52 ]	= 'hB6;
		virtual_vram[ 17'h07A53 ]	= 'hB8;
		virtual_vram[ 17'h07A54 ]	= 'hBC;
		virtual_vram[ 17'h07A55 ]	= 'hBC;
		virtual_vram[ 17'h07A56 ]	= 'hF8;
		virtual_vram[ 17'h07A57 ]	= 'h79;
		virtual_vram[ 17'h07A58 ]	= 'h79;
		virtual_vram[ 17'h07A59 ]	= 'h79;
		virtual_vram[ 17'h07A5A ]	= 'hF3;
		virtual_vram[ 17'h07A5B ]	= 'hF3;
		virtual_vram[ 17'h07A5C ]	= 'hFF;
		virtual_vram[ 17'h07A5D ]	= 'hDF;
		virtual_vram[ 17'h07A5E ]	= 'h3F;
		virtual_vram[ 17'h07A5F ]	= 'h3F;
		virtual_vram[ 17'h07A60 ]	= 'h2C;
		virtual_vram[ 17'h07A61 ]	= 'h1C;
		virtual_vram[ 17'h07A62 ]	= 'h18;
		virtual_vram[ 17'h07A63 ]	= 'h18;
		virtual_vram[ 17'h07A64 ]	= 'h18;
		virtual_vram[ 17'h07A65 ]	= 'h18;
		virtual_vram[ 17'h07A66 ]	= 'h18;
		virtual_vram[ 17'h07A67 ]	= 'h18;
		virtual_vram[ 17'h07A68 ]	= 'h30;
		virtual_vram[ 17'h07A69 ]	= 'h30;
		virtual_vram[ 17'h07A6A ]	= 'h30;
		virtual_vram[ 17'h07A6B ]	= 'h01;
		virtual_vram[ 17'h07A6C ]	= 'h01;
		virtual_vram[ 17'h07A6D ]	= 'h13;
		virtual_vram[ 17'h07A6E ]	= 'h0F;
		virtual_vram[ 17'h07A6F ]	= 'h1F;
		virtual_vram[ 17'h07A70 ]	= 'h21;
		virtual_vram[ 17'h07A71 ]	= 'h21;
		virtual_vram[ 17'h07A72 ]	= 'h49;
		virtual_vram[ 17'h07A73 ]	= 'h47;
		virtual_vram[ 17'h07A74 ]	= 'h43;
		virtual_vram[ 17'h07A75 ]	= 'h43;
		virtual_vram[ 17'h07A76 ]	= 'h07;
		virtual_vram[ 17'h07A77 ]	= 'h86;
		virtual_vram[ 17'h07A78 ]	= 'h86;
		virtual_vram[ 17'h07A79 ]	= 'h86;
		virtual_vram[ 17'h07A7A ]	= 'h0C;
		virtual_vram[ 17'h07A7B ]	= 'h0C;
		virtual_vram[ 17'h07A7C ]	= 'h00;
		virtual_vram[ 17'h07A7D ]	= 'h20;
		virtual_vram[ 17'h07A7E ]	= 'hC0;
		virtual_vram[ 17'h07A7F ]	= 'hC0;
		virtual_vram[ 17'h07A80 ]	= 'hB8;
		virtual_vram[ 17'h07A81 ]	= 'h78;
		virtual_vram[ 17'h07A82 ]	= 'h00;
		virtual_vram[ 17'h07A83 ]	= 'h00;
		virtual_vram[ 17'h07A84 ]	= 'h00;
		virtual_vram[ 17'h07A85 ]	= 'h00;
		virtual_vram[ 17'h07A86 ]	= 'h00;
		virtual_vram[ 17'h07A87 ]	= 'h00;
		virtual_vram[ 17'h07A88 ]	= 'h00;
		virtual_vram[ 17'h07A89 ]	= 'h00;
		virtual_vram[ 17'h07A8A ]	= 'h00;
		virtual_vram[ 17'h07A8B ]	= 'h00;
		virtual_vram[ 17'h07A8C ]	= 'h00;
		virtual_vram[ 17'h07A8D ]	= 'h00;
		virtual_vram[ 17'h07A8E ]	= 'h00;
		virtual_vram[ 17'h07A8F ]	= 'h00;
		virtual_vram[ 17'h07A90 ]	= 'h00;
		virtual_vram[ 17'h07A91 ]	= 'h00;
		virtual_vram[ 17'h07A92 ]	= 'h00;
		virtual_vram[ 17'h07A93 ]	= 'h00;
		virtual_vram[ 17'h07A94 ]	= 'h00;
		virtual_vram[ 17'h07A95 ]	= 'h00;
		virtual_vram[ 17'h07A96 ]	= 'h00;
		virtual_vram[ 17'h07A97 ]	= 'h00;
		virtual_vram[ 17'h07A98 ]	= 'h00;
		virtual_vram[ 17'h07A99 ]	= 'h00;
		virtual_vram[ 17'h07A9A ]	= 'h00;
		virtual_vram[ 17'h07A9B ]	= 'h00;
		virtual_vram[ 17'h07A9C ]	= 'h00;
		virtual_vram[ 17'h07A9D ]	= 'h00;
		virtual_vram[ 17'h07A9E ]	= 'h00;
		virtual_vram[ 17'h07A9F ]	= 'h00;
		virtual_vram[ 17'h07AA0 ]	= 'h47;
		virtual_vram[ 17'h07AA1 ]	= 'h87;
		virtual_vram[ 17'h07AA2 ]	= 'hFE;
		virtual_vram[ 17'h07AA3 ]	= 'h7C;
		virtual_vram[ 17'h07AA4 ]	= 'h00;
		virtual_vram[ 17'h07AA5 ]	= 'h00;
		virtual_vram[ 17'h07AA6 ]	= 'h00;
		virtual_vram[ 17'h07AA7 ]	= 'h00;
		virtual_vram[ 17'h07AA8 ]	= 'h00;
		virtual_vram[ 17'h07AA9 ]	= 'h00;
		virtual_vram[ 17'h07AAA ]	= 'h00;
		virtual_vram[ 17'h07AAB ]	= 'h00;
		virtual_vram[ 17'h07AAC ]	= 'h00;
		virtual_vram[ 17'h07AAD ]	= 'h00;
		virtual_vram[ 17'h07AAE ]	= 'h00;
		virtual_vram[ 17'h07AAF ]	= 'h00;
		virtual_vram[ 17'h07AB0 ]	= 'h3F;
		virtual_vram[ 17'h07AB1 ]	= 'h1F;
		virtual_vram[ 17'h07AB2 ]	= 'h00;
		virtual_vram[ 17'h07AB3 ]	= 'h00;
		virtual_vram[ 17'h07AB4 ]	= 'h00;
		virtual_vram[ 17'h07AB5 ]	= 'h00;
		virtual_vram[ 17'h07AB6 ]	= 'h00;
		virtual_vram[ 17'h07AB7 ]	= 'h00;
		virtual_vram[ 17'h07AB8 ]	= 'h00;
		virtual_vram[ 17'h07AB9 ]	= 'h00;
		virtual_vram[ 17'h07ABA ]	= 'h00;
		virtual_vram[ 17'h07ABB ]	= 'h00;
		virtual_vram[ 17'h07ABC ]	= 'h00;
		virtual_vram[ 17'h07ABD ]	= 'h00;
		virtual_vram[ 17'h07ABE ]	= 'h00;
		virtual_vram[ 17'h07ABF ]	= 'h00;
		virtual_vram[ 17'h07AC0 ]	= 'h00;
		virtual_vram[ 17'h07AC1 ]	= 'h00;
		virtual_vram[ 17'h07AC2 ]	= 'h00;
		virtual_vram[ 17'h07AC3 ]	= 'h00;
		virtual_vram[ 17'h07AC4 ]	= 'h00;
		virtual_vram[ 17'h07AC5 ]	= 'h00;
		virtual_vram[ 17'h07AC6 ]	= 'h00;
		virtual_vram[ 17'h07AC7 ]	= 'h00;
		virtual_vram[ 17'h07AC8 ]	= 'h00;
		virtual_vram[ 17'h07AC9 ]	= 'h00;
		virtual_vram[ 17'h07ACA ]	= 'h00;
		virtual_vram[ 17'h07ACB ]	= 'h00;
		virtual_vram[ 17'h07ACC ]	= 'h00;
		virtual_vram[ 17'h07ACD ]	= 'h00;
		virtual_vram[ 17'h07ACE ]	= 'h00;
		virtual_vram[ 17'h07ACF ]	= 'h00;

		repeat( 50 ) @( negedge CLK21M );
		RESET		= 0;
		repeat( 10 ) @( posedge CLK21M );

		repeat( 300000 ) begin
			BWINDOW_Y = (DOTCOUNTERYP >= 9'd0 && DOTCOUNTERYP <= 191 ) ? 1'b1 : 1'b0;
			REG_R1_SP_SIZE = 1'b1;
			REG_R1_SP_ZOOM = 1'b0;
			REG_R11R5_SP_ATR_ADDR = 'h01e00 >> 7;
			REG_R6_SP_GEN_ADDR = 'h03800 >> 11;
			REG_R8_COL0_ON = 1'b0;
			REG_R8_SP_OFF = 1'b0;
			REG_R23_VSTART_LINE = 8'd0;
			REG_R27_H_SCROLL = 3'd0;
			SPMODE2 = 1'b1;
			VRAMINTERLEAVEMODE = 1'b0;
			@( posedge CLK21M );
		end
		$finish;
	end
endmodule
